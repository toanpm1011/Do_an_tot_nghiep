`include "uvm.sv"
`include "uvm_macros.svh"
import  uvm_pkg::*;

`include "../src/aes_env/aes_interface.sv"

`include "../src/aes_agent/aes_transaction.sv"
`include "../src/aes_agent/aes_driver.sv"
`include "../src/aes_agent/aes_monitor.sv"
`include "../src/aes_agent/aes_sequencer.sv"
`include "../src/aes_agent/aes_sequence.sv"
`include "../src/aes_agent/aes_agent.sv"

`include "../src/aes_scoreboard/aes_scoreboard.sv"
`include "../src/aes_env/aes_env.sv"
`include "../src/aes_test/test.sv"
