// UVM TLM macros _decl: define 2 analysis import to connect to tx_agent and rx_agent
`uvm_analysis_imp_decl(_encrypt)
`uvm_analysis_imp_decl(_decrypt)

class aes_scoreboard extends uvm_scoreboard;  
	`uvm_component_utils(aes_scoreboard)

  uvm_analysis_imp_encrypt #(aes_encrypt_transaction, aes_scoreboard) encrypt_ap_imp;
  uvm_analysis_imp_decrypt #(aes_decrypt_transaction, aes_scoreboard) decrypt_ap_imp;
//-----------------------------------------------------------------------------
// function : new
//-----------------------------------------------------------------------------
  function new (string name = "aes_scoreboard", uvm_component parent = null);
    super.new (name, parent);
  endfunction : new 
//-----------------------------------------------------------------------------
// function : build_phase
//-----------------------------------------------------------------------------
  function void build_phase (uvm_phase phase);
    super.build_phase(phase);
    encrypt_ap_imp = new ("encrypt_ap_imp", this);
    decrypt_ap_imp = new ("decrypt_ap_imp", this);
  endfunction
//-----------------------------------------------------------------------------
// function : write_tx
// Compare data from TX_DUT
//-----------------------------------------------------------------------------
  virtual function void write_encrypt(aes_encrypt_transaction item);
  	//if (item.plain_text_in == item.plain_text_out) begin
      //`uvm_info ("UVM_INFO","ENCRYPT CHECK PASS!", UVM_LOW)
      ///$display("plain_text_in = %b , ", item.plain_text_in);//, item.plain_text_out); // plain_text_out = %b */
      //`uvm_error ("UVM_ERROR","CHECK Failed!")
  endfunction : write_encrypt
//-----------------------------------------------------------------------------
// function : write_rx
// Compare data from RX_DUT
//-----------------------------------------------------------------------------
  virtual function void write_decrypt(aes_decrypt_transaction item);
    // if (item.cipher_text_in == item.cipher_text_out) begin
       `uvm_info ("UVM_INFO","DECRYPT PASS!", UVM_LOW)
    //     $display("cipher_text_in = %b , cipher_text_out = %b", item.cipher_text_in, item.cipher_text_out);
    // end 
    // else 
    //   `uvm_error ("UVM_ERROR","RX Failed!")
	endfunction : write_decrypt

endclass : aes_scoreboard