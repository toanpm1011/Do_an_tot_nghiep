
`include "uvm.sv"
`include "uvm_macros.svh"
import  uvm_pkg::*;

`include "../src/aes_env/aes_interface.sv"

`include "../src/aes_encrypt/aes_encrypt_transaction.sv"
`include "../src/aes_encrypt/aes_encrypt_driver.sv"
`include "../src/aes_encrypt/aes_encrypt_monitor.sv"
`include "../src/aes_encrypt/aes_encrypt_sequencer.sv"
`include "../src/aes_encrypt/aes_encrypt_sequence.sv"
`include "../src/aes_encrypt/aes_encrypt_agent.sv"

`include "../src/aes_decrypt/aes_decrypt_transaction.sv"
`include "../src/aes_decrypt/aes_decrypt_driver.sv"
`include "../src/aes_decrypt/aes_decrypt_monitor.sv"
`include "../src/aes_decrypt/aes_decrypt_sequencer.sv"
`include "../src/aes_decrypt/aes_decrypt_sequence.sv"
`include "../src/aes_decrypt/aes_decrypt_agent.sv"

`include "../src/aes_env/aes_scoreboard.sv"
`include "../src/aes_env/aes_env.sv"
`include "../src/aes_test/test.sv"
