`include "uvm.sv"
`include "uvm_macros.svh"
import  uvm_pkg::*;

`include "../src/aes_env/aes_interface.sv"

`include "../src/aes_agent/aes_encrypt_transaction.sv"
`include "../src/aes_agent/aes_encrypt_driver.sv"
`include "../src/aes_agent/aes_encrypt_monitor.sv"
`include "../src/aes_agent/aes_encrypt_sequencer.sv"
`include "../src/aes_agent/aes_encrypt_sequence.sv"
`include "../src/aes_agent/aes_encrypt_agent.sv"

`include "../src/aes_scoreboard/aes_scoreboard.sv"
`include "../src/aes_env/aes_env.sv"
`include "../src/aes_test/test.sv"
