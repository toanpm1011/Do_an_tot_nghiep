// MixColumn function
//
`include "AES_Mul_func.sv"
